module break_addr(
output [15:0] addr
);

assign addr = 16'h444d;

endmodule
