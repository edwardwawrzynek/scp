module break_addr(
output [15:0] addr
);

assign addr = 15'hf270;

endmodule
